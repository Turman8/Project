// ECG分类器参数
parameter INPUT_DIM = 15;
parameter OUTPUT_DIM = 1;
parameter DATA_WIDTH = 16;
parameter FRAC_BITS = 8;
